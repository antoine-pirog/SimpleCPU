library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity microprogram_memory is
    port (
        addr : in  std_logic_vector(4 downto 0);
        data : out std_logic_vector(15 downto 0)
    );
end microprogram_memory;

architecture behavioral of microprogram_memory is
    type rom_array is array (0 to 31) of std_logic_vector(15 downto 0);
    constant rom_data : rom_array := (
        "00001" & '0' & "000" & "00010" & "00", -- @0x0000
        "00010" & '0' & "101" & "00000" & "10", -- @0x0001
        "00011" & '0' & "101" & "00001" & "10", -- @0x0002
        "00000" & '1' & "000" & "00000" & "00", -- @0x0003
        "00000" & '0' & "000" & "00000" & "00", -- @0x0004
        "00110" & '0' & "001" & "00000" & "11", -- @0x0005
        "00111" & '0' & "001" & "10000" & "11", -- @0x0006
        "00000" & '0' & "000" & "00000" & "00", -- @0x0007
        "01001" & '0' & "000" & "00000" & "00", -- @0x0008
        "01010" & '0' & "000" & "00100" & "00", -- @0x0009
        "00000" & '0' & "000" & "00000" & "00", -- @0x000A
        "01100" & '0' & "001" & "00010" & "01", -- @0x000B
        "01101" & '0' & "001" & "00001" & "01", -- @0x000C
        "00000" & '0' & "000" & "00000" & "00", -- @0x000D
        "01111" & '0' & "001" & "00010" & "01", -- @0x000E
        "10000" & '0' & "001" & "10000" & "01", -- @0x000F
        "10001" & '0' & "101" & "00000" & "10", -- @0x0010
        "10010" & '0' & "101" & "00001" & "10", -- @0x0011
        "00000" & '0' & "000" & "00000" & "00", -- @0x0012
        "10100" & '0' & "100" & "00000" & "00", -- @0x0013
        "10101" & '0' & "100" & "10000" & "00", -- @0x0014
        "00000" & '0' & "000" & "00000" & "00", -- @0x0015
        "10111" & '0' & "000" & "00000" & "00", -- @0x0016
        "11000" & '0' & "000" & "01000" & "00", -- @0x0017
        "00000" & '0' & "000" & "00000" & "00", -- @0x0018
        "11010" & '0' & "110" & "00000" & "00", -- @0x0019
        "11011" & '0' & "110" & "10000" & "00", -- @0x001A
        "00000" & '0' & "000" & "00000" & "00", -- @0x001B
        "11101" & '0' & "111" & "00000" & "00", -- @0x001C
        "11110" & '0' & "111" & "10000" & "00", -- @0x001D
        "00000" & '0' & "000" & "00000" & "00", -- @0x001E
        "11111" & '1' & "000" & "00000" & "00"  -- @0x001F
    );
begin
    data <= rom_data(to_integer(unsigned(addr)));
end architecture;